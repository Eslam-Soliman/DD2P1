*** SPICE deck for cell Sim{sch} from library tri-state_Inverter
*** Created on Fri Mar 29, 2019 15:33:48
*** Last revised on Sat Mar 30, 2019 14:18:45
*** Written on Sat Mar 30, 2019 14:18:45 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tri-state_Inverter__tri-state_inv1x4 FROM CELL tri-state_inv1x4{sch}
.SUBCKT tri-state_Inverter__tri-state_inv1x4 a c F _c
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F a net@80 gnd N L=0.2U W=1.2U
Mnmos@1 net@80 c gnd gnd N L=0.2U W=1.2U
Mnmos@2 gnd c net@80 gnd N L=0.2U W=1.2U
Mnmos@3 net@80 a F gnd N L=0.2U W=1.2U
Mpmos@0 net@69 a F vdd P L=0.2U W=3.5U
Mpmos@1 vdd _c net@69 vdd P L=0.2U W=3.5U
Mpmos@2 net@69 _c vdd vdd P L=0.2U W=3.5U
Mpmos@3 F a net@69 vdd P L=0.2U W=3.5U
.ENDS tri-state_Inverter__tri-state_inv1x4

.global gnd vdd

*** TOP LEVEL CELL: Sim{sch}
Xtri-stat@9 a vdd F gnd tri-state_Inverter__tri-state_inv1x4

* Spice Code nodes in cell cell 'Sim{sch}'
.step param factor LIST 1 2 4 8
*** SUBCIRCUIT first__INV1x1 FROM CELL first:INV1x1{sch}
.SUBCKT first__INV1x1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.2U W= {factor*0.3U}
Mpmos@0 vdd in out vdd P L=0.2U W= {factor*0.7U}
.ENDS first__INV1x1
Xinverter@2 F out2 first__INV1x1
.step param t LIST 0p 100p 400p 800p
Vdd vdd 0 DC 3.3
Vin1 a 0 pulse 0 3.3 5n {t/0.6 + 0.00000001f} {t/0.6 + 0.00000001f} 5n {10 + t/0.3}
.tran 0 15n
.measure tpdf
+ TRIG V(a) VAL= 1.65 RISE = 1
+ TARG V(F) VAL=1.65 FALL = 1
.measure tpdr
+ TRIG V(a) VAL = 1.65 FALL = 1
+ TARG V(F) VAL = 1.65 RISE = 1
.measure diff param = tpdr - tpdf
.include C:\Electric\scmos18.txt
.END
