*** SPICE deck for cell AOI22x2_sim{sch} from library AOI
*** Created on Fri Mar 29, 2019 17:42:12
*** Last revised on Sat Mar 30, 2019 15:21:20
*** Written on Sat Mar 30, 2019 15:21:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT AOI__AOI22x2 FROM CELL AOI22x2{sch}
.SUBCKT AOI__AOI22x2 F w x y z
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F y net@23 gnd N L=0.2U W=1.2U
Mnmos@1 net@23 x gnd gnd N L=0.2U W=1.2U
Mnmos@2 F z net@24 gnd N L=0.2U W=1.2U
Mnmos@3 net@24 w gnd gnd N L=0.2U W=1.2U
Mpmos@0 net@6 y F vdd P L=0.2U W=3.9U
Mpmos@1 vdd w net@6 vdd P L=0.2U W=3.9U
Mpmos@2 net@6 x F vdd P L=0.2U W=3.9U
Mpmos@3 vdd z net@6 vdd P L=0.2U W=3.9U
.ENDS AOI__AOI22x2

.global gnd vdd

*** TOP LEVEL CELL: AOI22x2_sim{sch}
XAOI22x2@0 F w x y z AOI__AOI22x2

* Spice Code nodes in cell cell 'AOI22x2_sim{sch}'
.step param p1 LIST 0 3.3
.step param p2 LIST 0 3.3
.step param p3 LIST 0 3.3
Vdd vdd 0 DC 3.3
Vin1 x 0 DC {p1}
Vin2 y 0 DC {p2}
Vin3 z 0 DC {p3}
Vin4 w 0 DC 0
.tran 0 15n
.measure tran OutputVoltage param v(F)
.include C:\Users\Dell\Desktop\scmos18.txt
.END
.END
