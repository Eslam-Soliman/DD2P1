*** SPICE deck for cell AOI22x1_sim{sch} from library AOI
*** Created on Fri Mar 29, 2019 17:00:17
*** Last revised on Fri Mar 29, 2019 17:07:39
*** Written on Fri Mar 29, 2019 17:52:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT AOI__AOI22x1 FROM CELL AOI22x1{sch}
.SUBCKT AOI__AOI22x1 f w x y z
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 f y net@0 gnd N L=0.2U W=0.6U
Mnmos@1 net@0 x gnd gnd N L=0.2U W=0.6U
Mnmos@2 f z net@1 gnd N L=0.2U W=0.6U
Mnmos@3 net@1 w gnd gnd N L=0.2U W=0.6U
Mpmos@0 net@23 y f vdd P L=0.2U W=2.1U
Mpmos@1 vdd w net@23 vdd P L=0.2U W=2.1U
Mpmos@2 net@23 x f vdd P L=0.2U W=2.1U
Mpmos@3 vdd z net@23 vdd P L=0.2U W=2.1U
.ENDS AOI__AOI22x1

.global gnd vdd

*** TOP LEVEL CELL: AOI22x1_sim{sch}
XAOI22x1@0 F w x y z AOI__AOI22x1

* Spice Code nodes in cell cell 'AOI22x1_sim{sch}'
.step param factor LIST 1 2 4 8
*** SUBCIRCUIT first__INV1x1 FROM CELL first:INV1x1{sch}
.SUBCKT first__INV1x1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.2U W= {factor*0.3U}
Mpmos@0 vdd in out vdd P L=0.2U W= {factor*0.7U}
.ENDS first__INV1x1
Xinverter@2 F out2 first__INV1x1
.step param t LIST 0p 100p 400p 800p
Vdd vdd 0 DC 3.3
Vin1 x 0 pulse 0 3.3 5n {t/0.6 + 0.00000001f} {t/0.6 + 0.00000001f} 5n {10 + t/0.3}
Vin2 y 0 DC 3.3
Vin3 z 0 DC 0
Vin4 w 0 DC 0
.tran 0 15n
.measure tpdf
+ TRIG V(x) VAL= 1.65 RISE = 1
+ TARG V(F) VAL=1.65 FALL = 1
.measure tpdr
+ TRIG V(x) VAL = 1.65 FALL = 1
+ TARG V(F) VAL = 1.65 RISE = 1
.measure diff param = tpdr - tpdf
.include C:\Electric\scmos18.txt
.END
