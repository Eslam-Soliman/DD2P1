*** SPICE deck for cell NAND2x1_sim{sch} from library NAND
*** Created on Thu Mar 28, 2019 10:56:29
*** Last revised on Sat Mar 30, 2019 14:54:54
*** Written on Sat Mar 30, 2019 14:54:56 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT NAND__NAND2x1 FROM CELL NAND2x1{sch}
.SUBCKT NAND__NAND2x1 a b F
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F b net@0 gnd N L=0.2U W=2.4U
Mnmos@1 net@0 a gnd gnd N L=0.2U W=2.4U
Mpmos@0 vdd b F vdd P L=0.2U W=4.2U
Mpmos@1 vdd a F vdd P L=0.2U W=4.2U
.ENDS NAND__NAND2x1

.global gnd vdd

*** TOP LEVEL CELL: NAND2x1_sim{sch}
XNAND2x1@0 a b F NAND__NAND2x1

* Spice Code nodes in cell cell 'NAND2x1_sim{sch}'
.step param p1 LIST 0 3.3
.step param p2 LIST 0 3.3
Vdd vdd 0 DC 3.3
Vin1 a 0 DC {p1}
Vin2 b 0 DC {p2}
.tran 0 15n
.measure tran OutputVoltage param v(F)
.include C:\Users\Dell\Desktop\scmos18.txt
.END
.END
