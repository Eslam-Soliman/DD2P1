*** SPICE deck for cell Sim{sch} from library NOR2
*** Created on Sat Mar 30, 2019 14:48:09
*** Last revised on Sat Mar 30, 2019 14:53:46
*** Written on Sat Mar 30, 2019 15:27:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT NOR2__NOR2x1 FROM CELL NOR2x1{sch}
.SUBCKT NOR2__NOR2x1 a b F gnd vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F a gnd gnd N L=0.2U W=0.3U
Mnmos@1 F b gnd gnd N L=0.2U W=0.3U
Mpmos@0 net@21 b F vdd P L=0.2U W=1U
Mpmos@1 vdd a net@21 vdd P L=0.2U W=1U
.ENDS NOR2__NOR2x1

.global gnd vdd

*** TOP LEVEL CELL: Sim{sch}
XNOR2x1@0 a gnd F gnd vdd NOR2__NOR2x1

* Spice Code nodes in cell cell 'Sim{sch}'
.step param factor LIST 1 2 4 8
*** SUBCIRCUIT first__INV1x1 FROM CELL first:INV1x1{sch}
.SUBCKT first__INV1x1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.2U W= {factor*0.3U}
Mpmos@0 vdd in out vdd P L=0.2U W= {factor*0.7U}
.ENDS first__INV1x1
Xinverter@2 F out2 first__INV1x1
.step param t LIST 0p 100p 400p 800p
Vdd vdd 0 DC 3.3
Vin1 a 0 pulse 0 3.3 5n {t/0.6 + 0.00000001f} {t/0.6 + 0.00000001f} 5n {10 + t/0.3}
.tran 0 15n
.measure tpdf
+ TRIG V(a) VAL= 1.65 RISE = 1
+ TARG V(F) VAL=1.65 FALL = 1
.measure tpdr
+ TRIG V(a) VAL = 1.65 FALL = 1
+ TARG V(F) VAL = 1.65 RISE = 1
.measure diff param = tpdr - tpdf
.include C:\Electric\scmos18.txt
.END
