*** SPICE deck for cell Sim{sch} from library tri-state_Inverter
*** Created on Fri Mar 29, 2019 15:33:48
*** Last revised on Sat Mar 30, 2019 17:07:47
*** Written on Sat Mar 30, 2019 17:07:48 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tri-state_Inverter__tri-state_inv1x4 FROM CELL tri-state_inv1x4{sch}
.SUBCKT tri-state_Inverter__tri-state_inv1x4 a c F _c
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F a net@80 gnd N L=0.2U W=1.2U
Mnmos@1 net@80 c gnd gnd N L=0.2U W=1.2U
Mnmos@2 gnd c net@80 gnd N L=0.2U W=1.2U
Mnmos@3 net@80 a F gnd N L=0.2U W=1.2U
Mpmos@0 net@69 a F vdd P L=0.2U W=3.5U
Mpmos@1 vdd _c net@69 vdd P L=0.2U W=3.5U
Mpmos@2 net@69 _c vdd vdd P L=0.2U W=3.5U
Mpmos@3 F a net@69 vdd P L=0.2U W=3.5U
.ENDS tri-state_Inverter__tri-state_inv1x4

.global gnd vdd

*** TOP LEVEL CELL: Sim{sch}
Xtri-stat@16 a c F i tri-state_Inverter__tri-state_inv1x4

* Spice Code nodes in cell cell 'Sim{sch}'
.step param p1 LIST 0 3.3
.step param p2 LIST 0 3.3
Vdd vdd 0 DC 3.3
Vin1 c 0 DC {p2}
Vin2 i 0 DC {3.3 - p2}
Vin3 a 0 DC {p1}
.tran 0 15n
.measure tran OutputVoltage param v(F)
.include C:\Electric\scmos18.txt
.END
.END
