*** SPICE deck for cell Sim{sch} from library tri-state_Inverter
*** Created on Fri Mar 29, 2019 15:33:48
*** Last revised on Fri Mar 29, 2019 16:08:32
*** Written on Fri Mar 29, 2019 16:08:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tri-state_Inverter__tri-state_inv1x1 FROM CELL tri-state_Inverter:tri-state_inv1x1{sch}
.SUBCKT tri-state_Inverter__tri-state_inv1x1 a c F _c
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F a net@3 gnd N L=0.2U W=0.6U
Mnmos@1 net@3 c gnd gnd N L=0.2U W=0.6U
Mpmos@0 net@1 a F vdd P L=0.2U W=1.4U
Mpmos@1 vdd _c net@1 vdd P L=0.2U W=1.4U
.ENDS tri-state_Inverter__tri-state_inv1x1

.global gnd vdd

*** TOP LEVEL CELL: tri-state_Inverter:Sim{sch}
Xtri-stat@0 tri-stat@0_a vdd tri-stat@0_F gnd tri-state_Inverter__tri-state_inv1x1

* Spice Code nodes in cell cell 'tri-state_Inverter:Sim{sch}'
Vdd vdd 0 DC 3.3
Vin1 a 0 pulse 0 3.3 5n {t/0.6 + 0.00000001f} {t/0.6 + 0.00000001f} 5n {10 + t/0.3}
.tran 0 15n
.measure tpdf
+ TRIG V(a) VAL= 1.65 RISE = 1
+ TARG V(F) VAL=1.65 FALL = 1
.measure tpdr
+ TRIG V(a) VAL = 1.65 FALL = 1
+ TARG V(F) VAL = 1.65 RISE = 1
.measure diff param = tpdr - tpdf
.include C:\Electric\scmos18.txt
.END
.END
