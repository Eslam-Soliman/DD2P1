*** SPICE deck for cell NAND2x4_sim{sch} from library NAND
*** Created on Fri Mar 29, 2019 15:56:27
*** Last revised on Fri Mar 29, 2019 16:35:03
*** Written on Fri Mar 29, 2019 16:47:48 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT NAND__NAND2x4 FROM CELL NAND2x4{sch}
.SUBCKT NAND__NAND2x4 a b F
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F b net@0 gnd N L=0.2U W=2.4U
Mnmos@1 net@0 a gnd gnd N L=0.2U W=2.4U
Mpmos@0 vdd b F vdd P L=0.2U W=2.9U
Mpmos@1 vdd a F vdd P L=0.2U W=2.9U
.ENDS NAND__NAND2x4

.global gnd vdd

*** TOP LEVEL CELL: NAND2x4_sim{sch}
XNAND2x4@0 a b F NAND__NAND2x4

* Spice Code nodes in cell cell 'NAND2x4_sim{sch}'
.step param factor LIST 1 2 4 8
*** SUBCIRCUIT first__INV1x1 FROM CELL first:INV1x1{sch}
.SUBCKT first__INV1x1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.2U W= {factor*0.3U}
Mpmos@0 vdd in out vdd P L=0.2U W= {factor*0.9U}
.ENDS first__INV1x1
Xinverter@2 F out2 first__INV1x1
.step param t LIST 0p 100p 400p 800p
Vdd vdd 0 DC 3.3
Vin1 a 0 DC 3.3
Vin3 b 0 pulse 0 3.3 5n {t/0.6 + 0.00000001f} {t/0.6 + 0.00000001f} 5n {10 + t/0.3}
.tran 0 15n
.measure tpdf
+ TRIG V(b) VAL= 1.65 RISE = 1
+ TARG V(F) VAL=1.65 FALL = 1
.measure tpdr
+ TRIG V(b) VAL = 1.65 FALL = 1
+ TARG V(F) VAL = 1.65 RISE = 1
.measure diff param = tpdr - tpdf
.include C:\Users\Dell\Desktop\scmos18.txt
.END
